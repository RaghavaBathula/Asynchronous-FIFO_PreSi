package my_pkg;

	`include "asyncf_transaction.sv"
	`include "asyncf_down_transaction.sv"
	
	`include "asyncf_up_sequencer.sv"
	`include "asyncf_down_sequencer.sv"
	
	`include "asyncf_up_seq.sv"
	`include "asyncf_down_seq.sv"
	
	`include "asyncf_virtual_sequencer.sv"
	
	`include "asyncf_driver.sv"
	`include "asyncf_down_driver.sv"
	
	`include "asyncf_up_monitor.sv"
	`include "asyncf_down_monitor.sv"
	
	`include "asyncf_up_agent.sv"
	`include "asyncf_down_agent.sv"
	
	`include "asyncf_model.sv"
	
	`include "coverage.sv"
	
	`include "asyncf_scoreboard.sv"
	
	`include "asyncf_env.sv"
	
	`include "asyncf_case0_seq.sv"
	
	`include "asyncf_case1_seq.sv"
	

endpackage: my_pkg