package pkg;
	int tx_count = 32;
	`include "transaction.sv"
	`include "generator.sv"
	`include "driver.sv"
	`include "env.sv"

endpackage: pkg